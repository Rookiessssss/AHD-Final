library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity shift32bit is
PORT(shiftlr: IN STD_LOGIC;
     din: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	  imm: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  dout: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
end shift32bit;

architecture Behavioral of shift32bit is
SIGNAL doutl,doutr: STD_LOGIC_VECTOR(31 DOWNTO 0);

begin

WITH shiftlr SELECT
dout<= doutl WHEN '0',
       doutr WHEN '1',
		 x"ffffffff" WHEN OTHERS;
		 
WITH imm(4 DOWNTO 0) SELECT
  doutl<= 
   din(30 DOWNTO 0) & din(31) WHEN "00001",
   din(29 DOWNTO 0) & din(31 DOWNTO 30) WHEN "00010",
   din(28 DOWNTO 0) & din(31 DOWNTO 29) WHEN "00011",
   din(27 DOWNTO 0) & din(31 DOWNTO 28) WHEN "00100",
	din(26 DOWNTO 0) & din(31 DOWNTO 27) WHEN "00101",
	din(25 DOWNTO 0) & din(31 DOWNTO 26) WHEN "00110",
	din(24 DOWNTO 0) & din(31 DOWNTO 25) WHEN "00111",
	din(23 DOWNTO 0) & din(31 DOWNTO 24) WHEN "01000",
	din(22 DOWNTO 0) & din(31 DOWNTO 23) WHEN "01001",
	din(21 DOWNTO 0) & din(31 DOWNTO 22) WHEN "01010",
	din(20 DOWNTO 0) & din(31 DOWNTO 21) WHEN "01011",
	din(19 DOWNTO 0) & din(31 DOWNTO 20) WHEN "01100",
	din(18 DOWNTO 0) & din(31 DOWNTO 19) WHEN "01101",
	din(17 DOWNTO 0) & din(31 DOWNTO 18) WHEN "01110",
	din(16 DOWNTO 0) & din(31 DOWNTO 17) WHEN "01111",
	din(15 DOWNTO 0) & din(31 DOWNTO 16) WHEN "10000",
	din(14 DOWNTO 0) & din(31 DOWNTO 15) WHEN "10001",
	din(13 DOWNTO 0) & din(31 DOWNTO 14) WHEN "10010",
	din(12 DOWNTO 0) & din(31 DOWNTO 13) WHEN "10011",
	din(11 DOWNTO 0) & din(31 DOWNTO 12) WHEN "10100",
	din(10 DOWNTO 0) & din(31 DOWNTO 11) WHEN "10101",
	din(9 DOWNTO 0) & din(31 DOWNTO 10) WHEN "10110",
	din(8 DOWNTO 0) & din(31 DOWNTO 9) WHEN "10111",
	din(7 DOWNTO 0) & din(31 DOWNTO 8) WHEN "11000",
	din(6 DOWNTO 0) & din(31 DOWNTO 7) WHEN "11001",
	din(5 DOWNTO 0) & din(31 DOWNTO 6) WHEN "11010",
	din(4 DOWNTO 0) & din(31 DOWNTO 5) WHEN "11011",
	din(3 DOWNTO 0) & din(31 DOWNTO 4) WHEN "11100",
   din(2 DOWNTO 0) & din(31 DOWNTO 3) WHEN "11101",
	din(1 DOWNTO 0) & din(31 DOWNTO 2) WHEN "11110",
	din(0) & din(31 DOWNTO 1)   WHEN "11111",
   din   WHEN OTHERS;

WITH imm(4 DOWNTO 0) SELECT
doutr<=	din( 0) & din(31 DOWNTO 1) WHEN "00001",
	din(1 DOWNTO 0) & din(31 DOWNTO 2) WHEN "00010",
	din(2 DOWNTO 0) & din(31 DOWNTO 3) WHEN "00011",
	din(3 DOWNTO 0) & din(31 DOWNTO 4) WHEN "00100",
	din(4 DOWNTO 0) & din(31 DOWNTO 5) WHEN "00101",
	din(5 DOWNTO 0) & din(31 DOWNTO 6) WHEN "00110",
	din(6 DOWNTO 0) & din(31 DOWNTO 7) WHEN "00111",
	din(7 DOWNTO 0) & din(31 DOWNTO 8) WHEN "01000",
	din(8 DOWNTO 0) & din(31 DOWNTO 9) WHEN "01001",
	din(9 DOWNTO 0) & din(31 DOWNTO 10) WHEN "01010",
	din(10 DOWNTO 0) & din(31 DOWNTO 11) WHEN "01011",
	din(11 DOWNTO 0) & din(31 DOWNTO 12) WHEN "01100",
	din(12 DOWNTO 0) & din(31 DOWNTO 13) WHEN "01101",
	din(13 DOWNTO 0) & din(31 DOWNTO 14) WHEN "01110",
	din(14 DOWNTO 0) & din(31 DOWNTO 15) WHEN "01111",
	din(15 DOWNTO 0) & din(31 DOWNTO 16) WHEN "10000",
	din(16 DOWNTO 0) & din(31 DOWNTO 17) WHEN "10001",
	din(17 DOWNTO 0) & din(31 DOWNTO 18) WHEN "10010",
	din(18 DOWNTO 0) & din(31 DOWNTO 19) WHEN "10011",
	din(19 DOWNTO 0) & din(31 DOWNTO 20) WHEN "10100",
	din(20 DOWNTO 0) & din(31 DOWNTO 21) WHEN "10101",
	din(21 DOWNTO 0) & din(31 DOWNTO 22) WHEN "10110",
	din(22 DOWNTO 0) & din(31 DOWNTO 23) WHEN "10111",
	din(23 DOWNTO 0) & din(31 DOWNTO 24) WHEN "11000",
	din(24 DOWNTO 0) & din(31 DOWNTO 25) WHEN "11001",
	din(25 DOWNTO 0) & din(31 DOWNTO 26) WHEN "11010",
	din(26 DOWNTO 0) & din(31 DOWNTO 27) WHEN "11011",
	din(27 DOWNTO 0) & din(31 DOWNTO 28) WHEN "11100",
	din(28 DOWNTO 0) & din(31 DOWNTO 29) WHEN "11101",
	din(29 DOWNTO 0) & din(31 DOWNTO 30) WHEN "11110",
	din(30 DOWNTO 0) & din( 31) WHEN "11111",
	din WHEN OTHERS;

end Behavioral;

